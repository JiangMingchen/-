LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ALU0 IS
PORT(
 AC, DR: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
 AIM: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
 ISUM: IN STD_LOGIC;
 ESUM: IN STD_LOGIC;
 ALU_OUT: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
 );
END ALU0;
ARCHITECTURE A OF ALU0 IS
SIGNAL ALU_TEMP: STD_LOGIC_VECTOR(15 DOWNTO 0):="0000000000000000";
SIGNAL BIT0,BIT1,BIT2,BIT3,BIT4,BIT5,BIT6,BIT7:STD_LOGIC_VECTOR(15 DOWNTO 0):="0000000000000000";
------------------------------------
-------------AIM指令----------------
--AIM="0001" -> ADD
--AIM="0010" -> SUB
--AIM="0011" -> AND
--AIM="0100" -> OR
--AIM="1101" -> MUL
------------------------------------

BEGIN
PROCESS(AIM,ISUM,ESUM,AC,DR)
 BEGIN
  IF(ISUM='1') THEN
   IF(AIM="0001") THEN ALU_TEMP<=AC+DR;
   ELSIF(AIM="0010") THEN ALU_TEMP<=AC-DR;
   ELSIF(AIM="0011") THEN ALU_TEMP<=AC AND DR;
   ELSIF(AIM="0100") THEN ALU_TEMP<=AC OR DR;
	ELSIF(AIM="1101") THEN
	IF(AC(0)='1') THEN BIT0<=("00000000" & DR(7 DOWNTO 0)); ELSE BIT0<="0000000000000000"; END IF;
	IF(AC(1)='1') THEN BIT1<=("0000000" & DR(7 DOWNTO 0) & '0'); ELSE BIT1<="0000000000000000"; END IF;
	IF(AC(2)='1') THEN BIT2<=("000000" & DR(7 DOWNTO 0) & "00"); ELSE BIT2<="0000000000000000"; END IF;
	IF(AC(3)='1') THEN BIT3<=("00000" & DR(7 DOWNTO 0) & "000"); ELSE BIT3<="0000000000000000"; END IF;
	IF(AC(4)='1') THEN BIT4<=("0000" & DR(7 DOWNTO 0) & "0000"); ELSE BIT4<="0000000000000000"; END IF;
	IF(AC(5)='1') THEN BIT5<=("000" & DR(7 DOWNTO 0) & "00000"); ELSE BIT5<="0000000000000000"; END IF;
	IF(AC(6)='1') THEN BIT6<=("00" & DR(7 DOWNTO 0) & "000000"); ELSE BIT6<="0000000000000000"; END IF;
	IF(AC(7)='1') THEN BIT7<=('0' & DR(7 DOWNTO 0) & "0000000"); ELSE BIT7<="0000000000000000"; END IF;
   END IF;
  END IF;
  IF(ESUM='1') THEN 
  IF(AIM="1101") THEN ALU_OUT<=(((BIT0+BIT1)+(BIT2+BIT3))+((BIT4+BIT5)+(BIT6+BIT7)));
  ELSE ALU_OUT<=ALU_TEMP; END IF;
  ELSE
   ALU_OUT<="ZZZZZZZZZZZZZZZZ";
  END IF;
END PROCESS;
END A; 