LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY ACC0 IS
PORT(
 ADATA_IN:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
 IA:IN STD_LOGIC;
 EA:IN STD_LOGIC;
 CLK:IN STD_LOGIC;
 ADATA_OUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
 );
END ACC0;
ARCHITECTURE A OF ACC0 IS
SIGNAL REGQ : STD_LOGIC_VECTOR(15 DOWNTO 0);
BEGIN
 PROCESS(CLK,IA,EA)
 BEGIN
 IF(CLK'EVENT AND CLK='1') THEN
 IF(IA='1') THEN
 REGQ<=ADATA_IN;
 END IF;
 END IF;
 END PROCESS;
 ADATA_OUT<=REGQ WHEN EA='1' ELSE "ZZZZZZZZZZZZZZZZ"; 
END A; 