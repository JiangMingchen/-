LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX0 IS
PORT(
 DATA0:IN STD_LOGIC_VECTOR(2 DOWNTO 0):="ZZZ";
 DATA1:IN STD_LOGIC_VECTOR(2 DOWNTO 0):="ZZZ";
 WR:IN STD_LOGIC:='0';
 CHOOSE:OUT STD_LOGIC_VECTOR(2 DOWNTO 0):="ZZZ"
 ); 
END MUX0;
ARCHITECTURE A OF MUX0 IS
--SIGNAL CHOOSE:STD_LOGIC_VECTOR(15 DOWNTO 0):="ZZZZZZZZZZZZZZZZ";
BEGIN
process(DATA0,DATA1,WR)
begin
if(WR='1') then
CHOOSE <= DATA1;
else
CHOOSE <= DATA0;
end if;
end process;
END A; 