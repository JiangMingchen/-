LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY RAM0 IS
 PORT(
 WR,CS:IN STD_LOGIC;
 DIN:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
 DOUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0):="0000000000000000";
 ADDR:IN STD_LOGIC_VECTOR(2 DOWNTO 0)
 );
END RAM0;
ARCHITECTURE A OF RAM0 IS
TYPE MEMORY IS ARRAY(0 TO 7) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
BEGIN
 PROCESS(CS,WR,ADDR)
 VARIABLE MEM: MEMORY;
 BEGIN
 IF (CS='0') THEN
 IF (WR='0') THEN
 MEM(CONV_INTEGER(ADDR(2 DOWNTO 0))):=DIN;
 ELSIF(WR='1') THEN
 DOUT <= MEM(CONV_INTEGER(ADDR(2 DOWNTO 0)));
 END IF;
 END IF;
 END PROCESS;
END A; 