LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DBUS0 IS
PORT(
 INDATA1:IN STD_LOGIC_VECTOR(15 DOWNTO 0):="ZZZZZZZZZZZZZZZZ";
 INDATA2:IN STD_LOGIC_VECTOR(15 DOWNTO 0):="ZZZZZZZZZZZZZZZZ";
 OUTDATA:OUT STD_LOGIC_VECTOR(15 DOWNTO 0):="ZZZZZZZZZZZZZZZZ"
 ); 
END DBUS0;
ARCHITECTURE A OF DBUS0 IS
SIGNAL TEMP:STD_LOGIC_VECTOR(15 DOWNTO 0);
BEGIN
PROCESS(INDATA1,INDATA2)
BEGIN
	IF NOT(INDATA2 = "ZZZZZZZZZZZZZZZZ") THEN
		TEMP <= INDATA2;
	ELSE
		TEMP <= INDATA1;
	END IF;
END PROCESS;
OUTDATA<=TEMP;
END A; 
